ENTITY SMANGA IS
	PORT( LIMIT_SMANGA : IN BIT;
	VERDE_SMANGA : OUT BIT;
	AMARELO_SMANGA : OUT BIT;
	VERMELHO_SMANGA : OUT BIT);
END SMANGA;

ARCHITECTURE CKT OF SMANGA IS

SIGNAL 

BEGIN
	
END CKT;
