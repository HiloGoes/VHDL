--ENB SEMPRE EM '1'
--SEMPRE DAR CLEAR ANTES
ENTITY CONTADOR_8 IS
	PORT( CLK_CONTADOR_8 : IN BIT;
	ENB_CONTADOR_8 : IN BIT;
	CLR_CONTADOR_8 : IN BIT;
	SAIDA_CONTADOR_8 : OUT BIT_VECTOR (7 DOWNTO 0)
	);
END CONTADOR_8;

ARCHITECTURE CKT OF CONTADOR_8 IS

SIGNAL QCLK : BIT_VECTOR(6 DOWNTO 0);
SIGNAL CLK_ENB_CONTADOR_8 : BIT;

COMPONENT FFJK IS
 port(clk,J,K,P,C:in bit;
   q,qb:out bit);
END COMPONENT;

BEGIN
  
CLK_ENB_CONTADOR_8 <= CLK_CONTADOR_8 AND ENB_CONTADOR_8;

BIT0: FFJK PORT MAP( 
	 J=>'1',
	 K=>'1',
	 clk=>CLK_ENB_CONTADOR_8,
	 P=>'1',
	 C=>CLR_CONTADOR_8,
	 q=>SAIDA_CONTADOR_8(0),
	 qb=>QCLK(0)
);
BIT1: FFJK PORT MAP( 
	 J=>'1',
	 K=>'1',
	 clk=>QCLK(0),
	 P=>'1',
	 C=>CLR_CONTADOR_8,
	 q=>SAIDA_CONTADOR_8(1),
	 qb=>QCLK(1)
);
BIT2: FFJK PORT MAP( 
	 J=>'1',
	 K=>'1',
	 CLK=>QCLK(1),
	 P=>'1',
	 C=>CLR_CONTADOR_8,
	 Q=>SAIDA_CONTADOR_8(2),
	 QB=>QCLK(2)
);
BIT3: FFJK PORT MAP( 
	 J=>'1',
	 K=>'1',
	 CLK=>QCLK(2),
	 P=>'1',
	 C=>CLR_CONTADOR_8,
	 Q=>SAIDA_CONTADOR_8(3),
	 QB=>QCLK(3)
);
BIT4: FFJK PORT MAP( 
	 J=>'1',
	 K=>'1',
	 CLK=>QCLK(3),
	 P=>'1',
	 C=>CLR_CONTADOR_8,
	 Q=>SAIDA_CONTADOR_8(4),
	 QB=>QCLK(4)
);
BIT5: FFJK PORT MAP( 
	 J=>'1',
	 K=>'1',
	 CLK=>QCLK(4),
	 P=>'1',
	 C=>CLR_CONTADOR_8,
	 Q=>SAIDA_CONTADOR_8(5),
	 QB=>QCLK(5)
);
BIT6: FFJK PORT MAP( 
	 J=>'1',
	 K=>'1',
	 CLK=>QCLK(5),
	 P=>'1',
	 C=>CLR_CONTADOR_8,
	 Q=>SAIDA_CONTADOR_8(6),
	 QB=>QCLK(6)
);
BIT7: FFJK PORT MAP( 
	 J=>'1',
	 K=>'1',
	 CLK=>QCLK(6),
	 P=>'1',
	 C=>CLR_CONTADOR_8,
	 Q=>SAIDA_CONTADOR_8(7)
);
END CKT;
