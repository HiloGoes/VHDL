ENTITY MUX IS
	PORT( ENTRADA : IN BIT_VECTOR (3 DOWNTO 0);
	SEL : IN BIT_VECTOR(1 DOWNTO 0);
	SAI : OUT BIT);
END MUX;

ARCHITECTURE CKT OF MUX IS

SIGNAL S1,S2,S3,S4 : BIT;

BEGIN
  S1<= (NOT SEL(0))AND(NOT SEL(1)) and ENTRADA(0);
  S2	<= (SEL(0))AND(NOT SEL(1)) and ENTRADA(1);
  S3 <= (NOT SEL(0))AND( SEL(1)) and ENTRADA(2);
  S4 <= (SEL(0))AND(SEL(1)) and ENTRADA(3);
 	SAI	<= S1 or S2 OR S3 OR S4;
END CKT;