ENTITY SCAJU IS
	PORT( LIMIT_SCAJU : IN BIT;
	VERDE_SCAJU : OUT BIT;
	AMARELO_SCAJU : OUT BIT;
	VERMELHO_SCAJU : OUT BIT);
END SCAJU;

ARCHITECTURE CKT OF SCAJU IS

SIGNAL 

BEGIN
	
END CKT;
