G /15/V   15
Y /5 /V   20 
V /15/G   35
V /5 /Y   40

M     C   S

G /25/V   25
Y /5 /V   30
V /5 /G   35
V /5 /Y   40

  